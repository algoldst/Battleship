`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Cal Poly SLO CPE 133
// Engineer: Darian Primer
// 
// Create Date: 11/20/2018 01:22:30 AM
// Design Name: Top file for Master basys board(player A).
//////////////////////////////////////////////////////////////////////////////////


module Slave_Top(
    input [15:0] A,
    input [15:0] B,
    input LDR1B,
    input LDR2B,
    input clr,
    input DispB,
    output LivB,
    output OKB,
    output [15:0] B_Attack,
    output [7:0] seg,
    output [3:0] an,
    output BTN1B,
    output BTN2B,
    output BTN3B
    );
    
    



endmodule